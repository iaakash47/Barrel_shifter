* /home/user/eSim-Workspace/Barrel_shifter/bareelshifter.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Mon Jan 31 16:56:06 2022

.lib "sky130_fd_pr/models/sky130.lib.spice" tt

* Sheet Name: /
xM16 Out_4 GND input_in3 GND sky130_fd_pr__nfet_01v8 
xM17 Out_4 GND input_in4 GND sky130_fd_pr__nfet_01v8 	
xM18 Out_4 GND input_in5 GND sky130_fd_pr__nfet_01v8 			
xM19 Out_4 GND input_in6 GND sky130_fd_pr__nfet_01v8 	  
xM20 Out_4 Vdd input_in7 GND sky130_fd_pr__nfet_01v8 	
xM11 Out_3 GND input_in2 GND sky130_fd_pr__nfet_01v8 		
xM12 Out_3 GND input_in3 GND sky130_fd_pr__nfet_01v8 		
xM13 Out_3 GND input_in4 GND sky130_fd_pr__nfet_01v8 		
xM14 Out_3 GND input_in5 GND sky130_fd_pr__nfet_01v8 	
xM15 Out_3 Vdd input_in6 GND sky130_fd_pr__nfet_01v8 		
xM6  Out_2 GND input_in1 GND sky130_fd_pr__nfet_01v8 		
xM7  Out_2 GND input_in2 GND sky130_fd_pr__nfet_01v8 
xM8  Out_2 GND input_in3 GND sky130_fd_pr__nfet_01v8 
xM9  Out_2 GND input_in4 GND sky130_fd_pr__nfet_01v8 
xM10 Out_2 Vdd input_in5 GND sky130_fd_pr__nfet_01v8		
xM1  Out_1 GND input_in0 GND sky130_fd_pr__nfet_01v8 	
xM2  Out_1 GND input_in1 GND sky130_fd_pr__nfet_01v8 			
xM3  Out_1 GND input_in2 GND sky130_fd_pr__nfet_01v8 		
xM4  Out_1 GND input_in3 GND sky130_fd_pr__nfet_01v8 	
xM5  Out_1 Vdd input_in4 GND sky130_fd_pr__nfet_01v8 			
*U1 input_in0 PORT
*U2 input_in1 PORT
*U3 input_in2 PORT
*U4 input_in3 PORT
*U5 Vdd PORT
*U6 input_in4 PORT
*U7 input_in5 PORT
*U8 input_in6 PORT
*U9 input_in7 PORT
*U10 Out_3 PORT
*U11 Out_2 PORT
*U12 Out_1 PORT
*U13 Out_4 PORT		

V1 input_in4 0 PULSE(0 1.8 1n 10p 10p 10n 20n)
V2 input_in5 0 PULSE(0 1.8 7n 10p 10p 10n 20n)
V3 input_in6 0 PULSE(0 1.8 3n 10p 10p 10n 20n)
V4 input_in7 0 PULSE(0 1.8 9n 10p 10p 10n 20n)
VDD Vdd 0 1.5V
V6 input_in0 0 PULSE(0 1.8 4n 10p 10p 10n 20n)
V7 input_in1 0 PULSE(0 1.8 8n 10p 10p 10n 20n)
V8 input_in2 0 PULSE(0 1.8 12n 10p 10p 10n 20n)
V9 input_in3 0 PULSE(0 1.8 16n 10p 10p 10n 20n)

.tran 0.4ns 40ns 

.control
run
plot V(input_in0)
plot V(input_in1) 
plot V(input_in2) 
plot V(input_in3) 
plot V(input_in4) 
plot V(input_in5) 
plot V(input_in6) 
plot V(input_in7)
plot V(Out_1)   
plot V(Out_2)
plot V(Out_3) 
plot V(Out_4)  


.endc
.end
